// Copyright (C) 2020 Intel Corporation.
// SPDX-License-Identifier: MIT

//
// Description
//-----------------------------------------------------------------------------
//
//   Top level testbench with OFS top level module instantiated as DUT
//
//-----------------------------------------------------------------------------

`include "vendor_defines.vh"
`include "fpga_defines.vh"

import ofs_fim_cfg_pkg::*;
import ofs_fim_if_pkg::*;
import ofs_fim_pcie_hdr_def::*;
import ofs_fim_pcie_pkg::*;
import ofs_fim_eth_if_pkg::*;
`ifdef INCLUDE_DDR4 
import ofs_fim_mem_if_pkg::*; 
`endif

task SOC_REQ_OFF;
begin
   force top_tb.DUT.soc_pcie_wrapper.pcie_top.tester.test_packet_sender.tx_packet = '{default:'0};
end
endtask

task SOC_REQ_ON;
begin
   release top_tb.DUT.soc_pcie_wrapper.pcie_top.tester.test_packet_sender.tx_packet;
end
endtask

task HOST_REQ_OFF;
begin
   force top_tb.DUT.pcie_wrapper.pcie_top.tester.test_packet_sender.tx_packet = '{default:'0};
end
endtask

task HOST_REQ_ON;
begin
   release top_tb.DUT.pcie_wrapper.pcie_top.tester.test_packet_sender.tx_packet;
end
endtask


module top_tb ();

logic SYS_REFCLK;
logic PCIE_REFCLK0;
logic PCIE_REFCLK1;
logic PCIE_RESET_N;
logic ETH_REFCLK;
logic flash_reset;

logic SOC_PCIE_REFCLK0;
logic SOC_PCIE_REFCLK1;
logic SOC_PCIE_RESET_N;
   
initial begin
   SYS_REFCLK   = 0;
   PCIE_REFCLK0 = 0;
   PCIE_REFCLK1 = 0;
   PCIE_RESET_N = 0;
   SOC_PCIE_REFCLK0 = 0;
   SOC_PCIE_REFCLK1 = 0;
   SOC_PCIE_RESET_N = 0;
   ETH_REFCLK   = 0;
   flash_reset  = 0;
`ifdef SIM_MODE_SOC
   HOST_REQ_OFF();
`else
   SOC_REQ_OFF();
`endif
end

initial 
begin
`ifdef VCD_ON  
   `ifndef VCD_OFF
        $vcdpluson;
        $vcdplusmemon();
   `endif 
`endif
end        

`ifdef INCLUDE_DDR4
   ofs_fim_emif_ddr4_if ddr4_mem     [ofs_fim_mem_if_pkg::NUM_MEM_CHANNELS-1:0] ();
`endif

`ifdef INCLUDE_HSSI
// HSSI serial data for loopback
ofs_fim_hssi_serial_if hssi_if [NUM_ETH_LANES-1:0]();
// CVL BFM serial port tx/rx wrt FPGA/DUT
logic [NUM_CVL_LANES-1:0] cvl_serial_tx_p;
logic [NUM_CVL_LANES-1:0] cvl_serial_rx_p;
`endif

`ifdef INCLUDE_PMCI                                                                              
  logic          qspi_dclk;                                                 
  logic          qspi_ncs;                                                  
  wire    [3:0]  qspi_data;
  wire           spi_ingress_sclk;  
  wire           spi_ingress_csn;   
  wire           spi_ingress_miso;  
  wire           spi_ingress_mosi;  
  wire           spi_egress_mosi;   
  wire           spi_egress_csn;    
  wire           spi_egress_sclk;   
  wire           spi_egress_miso;   
`endif

always #5000 SYS_REFCLK   = ~SYS_REFCLK;   // 100MHz

initial #2us SOC_PCIE_RESET_N = 1; //  IOPLL sim model requires at least 1us of reset
always #5000 SOC_PCIE_REFCLK0 = ~SOC_PCIE_REFCLK0; // 100MHz
always #5000 SOC_PCIE_REFCLK1 = ~SOC_PCIE_REFCLK1; // 100MHz
initial #2us PCIE_RESET_N = 1; //  IOPLL sim model requires at least 1us of reset
always #5000 PCIE_REFCLK0 = ~PCIE_REFCLK0; // 100MHz
always #5000 PCIE_REFCLK1 = ~PCIE_REFCLK1; // 100MHz
always #3200 ETH_REFCLK   = ~ETH_REFCLK;   // 156.25MHz
always #10000 flash_reset = 1;

top DUT (

 `ifdef INCLUDE_DDR4
   .ddr4_mem     (ddr4_mem),
 `endif 
 
 `ifdef INCLUDE_HSSI
    `ifdef PMCI_QSFP
       //to make QSFP connections without affecting HSSI operations
      .hssi_if          (hssi_if),
    `else
      .qsfp_ref_clk     (ETH_REFCLK),
      .hssi_if          (hssi_if),
    //`ifdef INCLUDE_CVL
    //.cvl_serial_tx_p  (cvl_serial_tx_p),
    //.cvl_serial_rx_p  (cvl_serial_rx_p),
    //`endif
 `endif
 `endif

`ifdef INCLUDE_PMCI                                                                              
  // AC FPGA - AC card BMC interface 
  .qspi_dclk (qspi_dclk),                                                 
  .qspi_ncs  (qspi_ncs),                                                  
  .qspi_data (qspi_data), 
`ifdef SPI_LB                                                                              
  .spi_ingress_sclk(spi_ingress_sclk),       
  .spi_ingress_csn(spi_ingress_csn),        
  .spi_ingress_miso(spi_ingress_miso),       
  .spi_ingress_mosi(spi_ingress_mosi),       
  .spi_egress_mosi(spi_ingress_mosi),        
  .spi_egress_csn(spi_ingress_csn),         
  .spi_egress_sclk(spi_ingress_sclk),        
  .spi_egress_miso(spi_ingress_miso),         
`endif 
`ifdef BMC_EN
  .spi_ingress_sclk(bmc_m10.ingr_spi_clk),       
  .spi_ingress_csn(bmc_m10.ingr_spi_csn),        
  .spi_ingress_miso(bmc_m10.ingr_spi_miso),       
  .spi_ingress_mosi(bmc_m10.ingr_spi_mosi),       
  .spi_egress_mosi(bmc_m10.egrs_spi_mosi),        
  .spi_egress_csn(bmc_m10.egrs_spi_csn),         
  .spi_egress_sclk(bmc_m10.egrs_spi_clk),        
  .spi_egress_miso(bmc_m10.egrs_spi_miso),         
`endif 
`endif  
 
   .SOC_PCIE_REFCLK0    (SOC_PCIE_REFCLK0),
   .SOC_PCIE_REFCLK1    (SOC_PCIE_REFCLK1),
   .SOC_PCIE_RESET_N    (SOC_PCIE_RESET_N),
   .SOC_PCIE_RX_P       ('0),
   .SOC_PCIE_RX_N       ('0),
   .SOC_PCIE_TX_P       (),
   .SOC_PCIE_TX_N       (),

  .SYS_REFCLK      (SYS_REFCLK),
  .PCIE_REFCLK0    (PCIE_REFCLK0),
  .PCIE_REFCLK1    (PCIE_REFCLK1),
  .PCIE_RESET_N    (PCIE_RESET_N),
  .PCIE_RX_P       ('0),
  .PCIE_RX_N       ('0),
  .PCIE_TX_P       (),
  .PCIE_TX_N       ()
);


`ifdef INCLUDE_PMCI                                                                              
// MT25QxxxTop DUT (S, C, HOLD_DQ3, DQ0, DQ1, Vcc, Vpp_W_DQ2, RESET2); 
   
/*   N25Qxxx N25Qxxx (.S (qspi_ncs), 
                    .C_ (qspi_dclk), 
               .HOLD_DQ3(qspi_data[3]),
               //.RESET_DQ3(qspi_data[3]), 
               .DQ0(qspi_data[0]), 
               .DQ1(qspi_data[1]), 
               .Vcc(1), 
               .Vpp_W_DQ2(qspi_data[2]));
*/

`ifdef BMC_EN
   bmc_top  bmc_m10 ();
`endif

`endif



// HSSI serial loopback
`ifdef INCLUDE_HSSI
  `ifdef PMCI_QSFP
  `else
      `ifdef LOOPBACK_CONNECTOR //looping same channel TX to RX
          assign hssi_if[0].rx_p = hssi_if[4].tx_p;
          assign hssi_if[1].rx_p = hssi_if[5].tx_p;
          assign hssi_if[2].rx_p = hssi_if[6].tx_p;
          assign hssi_if[3].rx_p = hssi_if[7].tx_p;
          assign hssi_if[4].rx_p = hssi_if[0].tx_p;
          assign hssi_if[5].rx_p = hssi_if[1].tx_p;
          assign hssi_if[6].rx_p = hssi_if[2].tx_p;
          assign hssi_if[7].rx_p = hssi_if[3].tx_p;
      `else
         `ifdef ETH_100G
             assign hssi_if[0].rx_p = hssi_if[4].tx_p;
             assign hssi_if[1].rx_p = hssi_if[5].tx_p;
             assign hssi_if[2].rx_p = hssi_if[6].tx_p;
             assign hssi_if[3].rx_p = hssi_if[7].tx_p;
             assign hssi_if[4].rx_p = hssi_if[0].tx_p;
             assign hssi_if[5].rx_p = hssi_if[1].tx_p;
             assign hssi_if[6].rx_p = hssi_if[2].tx_p;
             assign hssi_if[7].rx_p = hssi_if[3].tx_p;
         
        `else
             assign hssi_if[0].rx_p = hssi_if[1].tx_p;
             assign hssi_if[1].rx_p = hssi_if[2].tx_p;
             assign hssi_if[2].rx_p = hssi_if[3].tx_p;
             assign hssi_if[3].rx_p = hssi_if[4].tx_p;
             assign hssi_if[4].rx_p = hssi_if[5].tx_p;
             assign hssi_if[5].rx_p = hssi_if[6].tx_p;
             assign hssi_if[6].rx_p = hssi_if[7].tx_p;
             assign hssi_if[7].rx_p = hssi_if[0].tx_p;
         `endif                                                        
      `endif                                                        
   `endif
`endif

// EMIF memory model   
`ifdef INCLUDE_DDR4
   genvar ch;
   generate
      for(ch=0; ch < ofs_fim_mem_if_pkg::NUM_MEM_CHANNELS; ch = ch+1) begin : mem_model
         initial ddr4_mem[ch].ref_clk = '0;
         always #833 ddr4_mem[ch].ref_clk = ~ddr4_mem[ch].ref_clk; // 1200 MHz
         ed_sim_mem ddr_mem_inst (
            .mem_ck     (ddr4_mem[ch].ck),
            .mem_ck_n   (ddr4_mem[ch].ck_n),
            .mem_a      (ddr4_mem[ch].a),
            .mem_act_n  (ddr4_mem[ch].act_n),
            .mem_ba     (ddr4_mem[ch].ba),
            .mem_bg     (ddr4_mem[ch].bg),
            .mem_cke    (ddr4_mem[ch].cke),
            .mem_cs_n   (ddr4_mem[ch].cs_n),
            .mem_odt    (ddr4_mem[ch].odt),
            .mem_reset_n(ddr4_mem[ch].reset_n),
            .mem_par    (ddr4_mem[ch].par),
            .mem_alert_n(ddr4_mem[ch].alert_n),
            .mem_dqs    (ddr4_mem[ch].dqs),
            .mem_dqs_n  (ddr4_mem[ch].dqs_n),
            .mem_dq     (ddr4_mem[ch].dq),
            .mem_dbi_n  (ddr4_mem[ch].dbi_n)
         );
      end
   endgenerate
`endif

`ifdef INCLUDE_PMCI
  pmci_if  pmci_if_1();
`endif

   
endmodule
