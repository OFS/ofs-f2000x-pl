// Copyright (C) 2020 Intel Corporation.
// SPDX-License-Identifier: MIT

//
// Description
//-----------------------------------------------------------------------------
//
//  CSR address 
//
//-----------------------------------------------------------------------------
`ifndef __TEST_CSR_DEFS__
`define __TEST_CSR_DEFS__

package test_csr_defs;
   localparam PCIE_DFH           = 32'h0;
   localparam PCIE_SCRATCHPAD    = PCIE_DFH + 32'h8;
   localparam PCIE_STAT          = PCIE_DFH + 32'h10;
   localparam PCIE_UNUSED_OFFSET = PCIE_DFH + 32'hff8;
endpackage

`endif
