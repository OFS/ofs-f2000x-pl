// Copyright (C) 2021 Intel Corporation.
// SPDX-License-Identifier: MIT

//
// Description
//-----------------------------------------------------------------------------
//
// This package defines the parameters used in PF/VF Mux module
//
//-----------------------------------------------------------------------------
package top_cfg_pkg;
   import ofs_fim_cfg_pkg::*;

   // Parameters
   parameter NUM_HOST = 1;
   parameter NUM_PORT = 2;
 
   parameter  FIM_NUM_PF         = 2;
   parameter  FIM_NUM_VF         = 0;
   parameter  FIM_MAX_NUM_VF     = 0;
   parameter  FIM_PF_WIDTH       = (FIM_NUM_PF < 2) ? 1 : $clog2(FIM_NUM_PF);
   parameter  FIM_VF_WIDTH       = (FIM_NUM_VF < 2) ? 1 : $clog2(FIM_NUM_VF);
 
//-------------------------------------------------------------------
// PF/VF Mapping Table 
//
// Host AFU: 
//    +---------------------------------+
//    + Module          | PF/VF         +
//    +---------------------------------+
//    | ST2MM           | PF0           | 
//    | HE-LB           | PF1           |
//    +---------------------------------+
//
//
//-------------------------------------------------------------------
//------------------------------------------------------------------------------------------------------------------------------------------------------
//  Physical Function#       Virtual Active           Virtual Function#        Switch/Mux Port ID        // AXI-S Pipeline Depth        // FPGA Device PF/VF to Switch Port Map
//------------------------------------------------------------------------------------------------------------------------------------------------------

   // ----- Mapping Table Begin -----
   // PF/VF Port IDs
   parameter SR_PF0_PF0_PID = 0;
   parameter SR_PF1_PF1_PID = 1;
  
   //=========================================================================================================================
   //                           PF/VF Mux Routing Table
   //=========================================================================================================================

   // The routing table is passed to the main PF/VF MUX instantiated in afu_top.
   // The PF/VF MUX has a function that parses the table in order to generate
   // a routing network.

   // Routing Table
   localparam NUM_RTABLE_ENTRIES = NUM_PORT+2;
    
   parameter NID_WIDTH = $clog2(NUM_PORT);// ID field width for targeting mux ports
   parameter MID_WIDTH = $clog2(NUM_HOST);// ID field width for targeting host ports
  
   // Number of MUX ports connected to the static region
   localparam NUM_SR_PORTS = NUM_PORT;

   // PF/VF mapping for FIM AFUs
   localparam int          AFU_SR_MUX_PID        [NUM_SR_PORTS] = '{SR_PF0_PF0_PID, SR_PF1_PF1_PID};
   localparam logic [11:0] PG_SR_PORTS_VF_NUM    [NUM_SR_PORTS] = '{0, 0}; 
   localparam logic        PG_SR_PORTS_VF_ACTIVE [NUM_SR_PORTS] = '{0, 0}; 
   localparam logic [2:0]  PG_SR_PORTS_PF_NUM    [NUM_SR_PORTS] = '{0, 1}; 

   
   import pcie_ss_hdr_pkg::ReqHdr_pf_vf_info_t;
   typedef pcie_ss_hdr_pkg::ReqHdr_pf_vf_info_t [NUM_SR_PORTS-1:0] t_sr_afu_pf_vf_info;
   typedef pf_vf_mux_pkg::t_pfvf_rtable_entry [NUM_RTABLE_ENTRIES-1:0] t_pf_vf_entry_info;

   function automatic t_sr_afu_pf_vf_info get_sr_pf_vf_info();
      t_sr_afu_pf_vf_info map;
      for (int p = 0; p < NUM_SR_PORTS; p = p + 1) begin
	 map[p].pf_num    = PG_SR_PORTS_PF_NUM[p];
	 map[p].vf_num    = PG_SR_PORTS_VF_NUM[p];
	 map[p].vf_active = PG_SR_PORTS_VF_ACTIVE[p];
      end
      return map;
   endfunction // gen_pf_vf_map

   // Sets the routing table in Static Region
   // Sets the PID routing information in fim_afu_instances
    function automatic t_pf_vf_entry_info get_pf_vf_entry_info();
      t_pf_vf_entry_info map;
      for (int p = 0; p < NUM_RTABLE_ENTRIES; p = p + 1) begin
         if(p<NUM_SR_PORTS) begin                        // Updates the routing table entry for all functions
            map[p].pf        = PG_SR_PORTS_PF_NUM[p];       // in the static region
	    map[p].vf        = PG_SR_PORTS_VF_NUM[p];
	    map[p].vf_active = PG_SR_PORTS_VF_ACTIVE[p];
            map[p].pfvf_port = AFU_SR_MUX_PID[p];
         end else begin                                     //Default entries that are mapped to PID 0 always
            map[p].pf    = -1;
	    map[p].vf    = -1;
	    map[p].vf_active = (p == (NUM_RTABLE_ENTRIES-1));
            map[p].pfvf_port = 0;
         end
      end
      return map;
   endfunction // gen_pf_vf_map

endpackage : top_cfg_pkg
