// Copyright (C) 2022 Intel Corporation.
// SPDX-License-Identifier: MIT

// Description
//-----------------------------------------------------------------------------
// Host AFU Peripheral Fabric interface wrapper
//-----------------------------------------------------------------------------

module apf_top (
   input logic clk,
   input logic rst_n,

   // APF managers
   ofs_fim_axi_lite_if.slave apf_st2mm_mst_if,
   ofs_fim_axi_lite_if.slave apf_bpf_mst_if,
   ofs_fim_axi_lite_if.slave apf_mctp_mst_if, 
   // APF functions
   ofs_fim_axi_lite_if.master apf_achk_slv_if,
   ofs_fim_axi_lite_if.master apf_bpf_slv_if,
   ofs_fim_axi_lite_if.master apf_st2mm_slv_if
);
		
  apf apf_inst (
   .clk_clk             (clk),
   .rst_n_reset_n       (rst_n),

   .apf_bpf_mst_awaddr  (apf_bpf_mst_if.awaddr),
   .apf_bpf_mst_awprot  (apf_bpf_mst_if.awprot),
   .apf_bpf_mst_awvalid (apf_bpf_mst_if.awvalid),
   .apf_bpf_mst_awready (apf_bpf_mst_if.awready),
   .apf_bpf_mst_wdata   (apf_bpf_mst_if.wdata),
   .apf_bpf_mst_wstrb   (apf_bpf_mst_if.wstrb),
   .apf_bpf_mst_wvalid  (apf_bpf_mst_if.wvalid),
   .apf_bpf_mst_wready  (apf_bpf_mst_if.wready),
   .apf_bpf_mst_bresp   (apf_bpf_mst_if.bresp),
   .apf_bpf_mst_bvalid  (apf_bpf_mst_if.bvalid),
   .apf_bpf_mst_bready  (apf_bpf_mst_if.bready),
   .apf_bpf_mst_araddr  (apf_bpf_mst_if.araddr),
   .apf_bpf_mst_arprot  (apf_bpf_mst_if.arprot),
   .apf_bpf_mst_arvalid (apf_bpf_mst_if.arvalid),
   .apf_bpf_mst_arready (apf_bpf_mst_if.arready),
   .apf_bpf_mst_rdata   (apf_bpf_mst_if.rdata),
   .apf_bpf_mst_rresp   (apf_bpf_mst_if.rresp),
   .apf_bpf_mst_rvalid  (apf_bpf_mst_if.rvalid),
   .apf_bpf_mst_rready  (apf_bpf_mst_if.rready),

   .apf_st2mm_mst_awaddr  ( apf_st2mm_mst_if.awaddr),
   .apf_st2mm_mst_awprot  ( apf_st2mm_mst_if.awprot),
   .apf_st2mm_mst_awvalid ( apf_st2mm_mst_if.awvalid),
   .apf_st2mm_mst_awready ( apf_st2mm_mst_if.awready),
   .apf_st2mm_mst_wdata   ( apf_st2mm_mst_if.wdata),
   .apf_st2mm_mst_wstrb   ( apf_st2mm_mst_if.wstrb),
   .apf_st2mm_mst_wvalid  ( apf_st2mm_mst_if.wvalid),
   .apf_st2mm_mst_wready  ( apf_st2mm_mst_if.wready),
   .apf_st2mm_mst_bresp   ( apf_st2mm_mst_if.bresp),
   .apf_st2mm_mst_bvalid  ( apf_st2mm_mst_if.bvalid),
   .apf_st2mm_mst_bready  ( apf_st2mm_mst_if.bready),
   .apf_st2mm_mst_araddr  ( apf_st2mm_mst_if.araddr),
   .apf_st2mm_mst_arprot  ( apf_st2mm_mst_if.arprot),
   .apf_st2mm_mst_arvalid ( apf_st2mm_mst_if.arvalid),
   .apf_st2mm_mst_arready ( apf_st2mm_mst_if.arready),
   .apf_st2mm_mst_rdata   ( apf_st2mm_mst_if.rdata),
   .apf_st2mm_mst_rresp   ( apf_st2mm_mst_if.rresp),
   .apf_st2mm_mst_rvalid  ( apf_st2mm_mst_if.rvalid),
   .apf_st2mm_mst_rready  ( apf_st2mm_mst_if.rready),

   .apf_mctp_mst_awaddr  ( apf_mctp_mst_if.awaddr),
   .apf_mctp_mst_awprot  ( apf_mctp_mst_if.awprot),
   .apf_mctp_mst_awvalid ( apf_mctp_mst_if.awvalid),
   .apf_mctp_mst_awready ( apf_mctp_mst_if.awready),
   .apf_mctp_mst_wdata   ( apf_mctp_mst_if.wdata),
   .apf_mctp_mst_wstrb   ( apf_mctp_mst_if.wstrb),
   .apf_mctp_mst_wvalid  ( apf_mctp_mst_if.wvalid),
   .apf_mctp_mst_wready  ( apf_mctp_mst_if.wready),
   .apf_mctp_mst_bresp   ( apf_mctp_mst_if.bresp),
   .apf_mctp_mst_bvalid  ( apf_mctp_mst_if.bvalid),
   .apf_mctp_mst_bready  ( apf_mctp_mst_if.bready),
   .apf_mctp_mst_araddr  ( apf_mctp_mst_if.araddr),
   .apf_mctp_mst_arprot  ( apf_mctp_mst_if.arprot),
   .apf_mctp_mst_arvalid ( apf_mctp_mst_if.arvalid),
   .apf_mctp_mst_arready ( apf_mctp_mst_if.arready),
   .apf_mctp_mst_rdata   ( apf_mctp_mst_if.rdata),
   .apf_mctp_mst_rresp   ( apf_mctp_mst_if.rresp),
   .apf_mctp_mst_rvalid  ( apf_mctp_mst_if.rvalid),
   .apf_mctp_mst_rready  ( apf_mctp_mst_if.rready),
   
   .apf_achk_slv_awaddr  (apf_achk_slv_if.awaddr),
   .apf_achk_slv_awprot  (apf_achk_slv_if.awprot),
   .apf_achk_slv_awvalid (apf_achk_slv_if.awvalid),
   .apf_achk_slv_awready (apf_achk_slv_if.awready),
   .apf_achk_slv_wdata   (apf_achk_slv_if.wdata),
   .apf_achk_slv_wstrb   (apf_achk_slv_if.wstrb),
   .apf_achk_slv_wvalid  (apf_achk_slv_if.wvalid),
   .apf_achk_slv_wready  (apf_achk_slv_if.wready),
   .apf_achk_slv_bresp   (apf_achk_slv_if.bresp),
   .apf_achk_slv_bvalid  (apf_achk_slv_if.bvalid),
   .apf_achk_slv_bready  (apf_achk_slv_if.bready),
   .apf_achk_slv_araddr  (apf_achk_slv_if.araddr),
   .apf_achk_slv_arprot  (apf_achk_slv_if.arprot),
   .apf_achk_slv_arvalid (apf_achk_slv_if.arvalid),
   .apf_achk_slv_arready (apf_achk_slv_if.arready),
   .apf_achk_slv_rdata   (apf_achk_slv_if.rdata),
   .apf_achk_slv_rresp   (apf_achk_slv_if.rresp),
   .apf_achk_slv_rvalid  (apf_achk_slv_if.rvalid),
   .apf_achk_slv_rready  (apf_achk_slv_if.rready),
 
   .apf_bpf_slv_awaddr  (apf_bpf_slv_if.awaddr),
   .apf_bpf_slv_awprot  (apf_bpf_slv_if.awprot),
   .apf_bpf_slv_awvalid (apf_bpf_slv_if.awvalid),
   .apf_bpf_slv_awready (apf_bpf_slv_if.awready),
   .apf_bpf_slv_wdata   (apf_bpf_slv_if.wdata),
   .apf_bpf_slv_wstrb   (apf_bpf_slv_if.wstrb),
   .apf_bpf_slv_wvalid  (apf_bpf_slv_if.wvalid),
   .apf_bpf_slv_wready  (apf_bpf_slv_if.wready),
   .apf_bpf_slv_bresp   (apf_bpf_slv_if.bresp),
   .apf_bpf_slv_bvalid  (apf_bpf_slv_if.bvalid),
   .apf_bpf_slv_bready  (apf_bpf_slv_if.bready),
   .apf_bpf_slv_araddr  (apf_bpf_slv_if.araddr),
   .apf_bpf_slv_arprot  (apf_bpf_slv_if.arprot),
   .apf_bpf_slv_arvalid (apf_bpf_slv_if.arvalid),
   .apf_bpf_slv_arready (apf_bpf_slv_if.arready),
   .apf_bpf_slv_rdata   (apf_bpf_slv_if.rdata),
   .apf_bpf_slv_rresp   (apf_bpf_slv_if.rresp),
   .apf_bpf_slv_rvalid  (apf_bpf_slv_if.rvalid),
   .apf_bpf_slv_rready  (apf_bpf_slv_if.rready),

   .apf_st2mm_slv_awaddr  ( apf_st2mm_slv_if.awaddr),
   .apf_st2mm_slv_awprot  ( apf_st2mm_slv_if.awprot),
   .apf_st2mm_slv_awvalid ( apf_st2mm_slv_if.awvalid),
   .apf_st2mm_slv_awready ( apf_st2mm_slv_if.awready),
   .apf_st2mm_slv_wdata   ( apf_st2mm_slv_if.wdata),
   .apf_st2mm_slv_wstrb   ( apf_st2mm_slv_if.wstrb),
   .apf_st2mm_slv_wvalid  ( apf_st2mm_slv_if.wvalid),
   .apf_st2mm_slv_wready  ( apf_st2mm_slv_if.wready),
   .apf_st2mm_slv_bresp   ( apf_st2mm_slv_if.bresp),
   .apf_st2mm_slv_bvalid  ( apf_st2mm_slv_if.bvalid),
   .apf_st2mm_slv_bready  ( apf_st2mm_slv_if.bready),
   .apf_st2mm_slv_araddr  ( apf_st2mm_slv_if.araddr),
   .apf_st2mm_slv_arprot  ( apf_st2mm_slv_if.arprot),
   .apf_st2mm_slv_arvalid ( apf_st2mm_slv_if.arvalid),
   .apf_st2mm_slv_arready ( apf_st2mm_slv_if.arready),
   .apf_st2mm_slv_rdata   ( apf_st2mm_slv_if.rdata),
   .apf_st2mm_slv_rresp   ( apf_st2mm_slv_if.rresp),
   .apf_st2mm_slv_rvalid  ( apf_st2mm_slv_if.rvalid),
   .apf_st2mm_slv_rready  ( apf_st2mm_slv_if.rready)

   );

endmodule
