// Copyright (C) 2023 Intel Corporation
// SPDX-License-Identifier: MIT

`ifndef TEST_TOP_PKG_SVH
`define TEST_TOP_PKG_SVH

    `include "test_pkg.svh"
    `include "test_long_pkg.svh"


`endif // TEST_TOP_PKG_SVH
