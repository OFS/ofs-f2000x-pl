// Copyright (C) 2022 Intel Corporation.
// SPDX-License-Identifier: MIT

// Description
//-----------------------------------------------------------------------------
// Board Peripheral Fabric interface wrapper
//-----------------------------------------------------------------------------

module bpf_top (
   input logic clk,
   input logic rst_n,

   // BPF managers
   ofs_fim_axi_lite_if.slave bpf_host_apf_mst_if,
   ofs_fim_axi_lite_if.slave bpf_soc_apf_mst_if,
   ofs_fim_axi_lite_if.slave bpf_fme_mst_if,
   ofs_fim_axi_lite_if.slave bpf_pmci_mst_if,
   // BPF functions
   ofs_fim_axi_lite_if.master bpf_pcie_slv_if,
   ofs_fim_axi_lite_if.master bpf_fme_slv_if,
   ofs_fim_axi_lite_if.master bpf_soc_apf_slv_if,
   ofs_fim_axi_lite_if.master bpf_soc_pcie_slv_if,
   ofs_fim_axi_lite_if.master bpf_emif_slv_if,
   ofs_fim_axi_lite_if.master bpf_hssi_slv_if,
   ofs_fim_axi_lite_if.master bpf_qsfp0_slv_if,
   ofs_fim_axi_lite_if.master bpf_qsfp1_slv_if,
   ofs_fim_axi_lite_if.master bpf_host_apf_slv_if,
   ofs_fim_axi_lite_if.master bpf_pmci_slv_if

);


bpf 
bpf_inst (
   .clk_clk                   (clk                       ),
   .rst_n_reset_n             (rst_n                     ),
   
   .bpf_apf_mst_awaddr        (bpf_soc_apf_mst_if.awaddr     ),
   .bpf_apf_mst_awprot        (bpf_soc_apf_mst_if.awprot     ),
   .bpf_apf_mst_awvalid       (bpf_soc_apf_mst_if.awvalid    ),
   .bpf_apf_mst_awready       (bpf_soc_apf_mst_if.awready    ),
   .bpf_apf_mst_wdata         (bpf_soc_apf_mst_if.wdata      ),
   .bpf_apf_mst_wstrb         (bpf_soc_apf_mst_if.wstrb      ),
   .bpf_apf_mst_wvalid        (bpf_soc_apf_mst_if.wvalid     ),
   .bpf_apf_mst_wready        (bpf_soc_apf_mst_if.wready     ),
   .bpf_apf_mst_bresp         (bpf_soc_apf_mst_if.bresp      ),
   .bpf_apf_mst_bvalid        (bpf_soc_apf_mst_if.bvalid     ),
   .bpf_apf_mst_bready        (bpf_soc_apf_mst_if.bready     ),
   .bpf_apf_mst_araddr        (bpf_soc_apf_mst_if.araddr     ),
   .bpf_apf_mst_arprot        (bpf_soc_apf_mst_if.arprot     ),
   .bpf_apf_mst_arvalid       (bpf_soc_apf_mst_if.arvalid    ),
   .bpf_apf_mst_arready       (bpf_soc_apf_mst_if.arready    ),
   .bpf_apf_mst_rdata         (bpf_soc_apf_mst_if.rdata      ),
   .bpf_apf_mst_rresp         (bpf_soc_apf_mst_if.rresp      ),
   .bpf_apf_mst_rvalid        (bpf_soc_apf_mst_if.rvalid     ),
   .bpf_apf_mst_rready        (bpf_soc_apf_mst_if.rready     ),
   
   .bpf_host_apf_mst_awaddr   (bpf_host_apf_mst_if.awaddr     ),
   .bpf_host_apf_mst_awprot   (bpf_host_apf_mst_if.awprot     ),
   .bpf_host_apf_mst_awvalid  (bpf_host_apf_mst_if.awvalid    ),
   .bpf_host_apf_mst_awready  (bpf_host_apf_mst_if.awready    ),
   .bpf_host_apf_mst_wdata    (bpf_host_apf_mst_if.wdata      ),
   .bpf_host_apf_mst_wstrb    (bpf_host_apf_mst_if.wstrb      ),
   .bpf_host_apf_mst_wvalid   (bpf_host_apf_mst_if.wvalid     ),
   .bpf_host_apf_mst_wready   (bpf_host_apf_mst_if.wready     ),
   .bpf_host_apf_mst_bresp    (bpf_host_apf_mst_if.bresp      ),
   .bpf_host_apf_mst_bvalid   (bpf_host_apf_mst_if.bvalid     ),
   .bpf_host_apf_mst_bready   (bpf_host_apf_mst_if.bready     ),
   .bpf_host_apf_mst_araddr   (bpf_host_apf_mst_if.araddr     ),
   .bpf_host_apf_mst_arprot   (bpf_host_apf_mst_if.arprot     ),
   .bpf_host_apf_mst_arvalid  (bpf_host_apf_mst_if.arvalid    ),
   .bpf_host_apf_mst_arready  (bpf_host_apf_mst_if.arready    ),
   .bpf_host_apf_mst_rdata    (bpf_host_apf_mst_if.rdata      ),
   .bpf_host_apf_mst_rresp    (bpf_host_apf_mst_if.rresp      ),
   .bpf_host_apf_mst_rvalid   (bpf_host_apf_mst_if.rvalid     ),
   .bpf_host_apf_mst_rready   (bpf_host_apf_mst_if.rready     ),
         
   .bpf_pcie_slv_awaddr       (bpf_pcie_slv_if.awaddr    ), 
   .bpf_pcie_slv_awprot       (bpf_pcie_slv_if.awprot    ), 
   .bpf_pcie_slv_awvalid      (bpf_pcie_slv_if.awvalid   ), 
   .bpf_pcie_slv_awready      (bpf_pcie_slv_if.awready   ), 
   .bpf_pcie_slv_wdata        (bpf_pcie_slv_if.wdata     ), 
   .bpf_pcie_slv_wstrb        (bpf_pcie_slv_if.wstrb     ), 
   .bpf_pcie_slv_wvalid       (bpf_pcie_slv_if.wvalid    ), 
   .bpf_pcie_slv_wready       (bpf_pcie_slv_if.wready    ), 
   .bpf_pcie_slv_bresp        (bpf_pcie_slv_if.bresp     ), 
   .bpf_pcie_slv_bvalid       (bpf_pcie_slv_if.bvalid    ), 
   .bpf_pcie_slv_bready       (bpf_pcie_slv_if.bready    ), 
   .bpf_pcie_slv_araddr       (bpf_pcie_slv_if.araddr    ), 
   .bpf_pcie_slv_arprot       (bpf_pcie_slv_if.arprot    ), 
   .bpf_pcie_slv_arvalid      (bpf_pcie_slv_if.arvalid   ), 
   .bpf_pcie_slv_arready      (bpf_pcie_slv_if.arready   ), 
   .bpf_pcie_slv_rdata        (bpf_pcie_slv_if.rdata     ), 
   .bpf_pcie_slv_rresp        (bpf_pcie_slv_if.rresp     ), 
   .bpf_pcie_slv_rvalid       (bpf_pcie_slv_if.rvalid    ), 
   .bpf_pcie_slv_rready       (bpf_pcie_slv_if.rready    ),

   .bpf_soc_pcie_slv_awaddr    (bpf_soc_pcie_slv_if.awaddr    ), 
   .bpf_soc_pcie_slv_awprot    (bpf_soc_pcie_slv_if.awprot    ), 
   .bpf_soc_pcie_slv_awvalid   (bpf_soc_pcie_slv_if.awvalid   ), 
   .bpf_soc_pcie_slv_awready   (bpf_soc_pcie_slv_if.awready   ), 
   .bpf_soc_pcie_slv_wdata     (bpf_soc_pcie_slv_if.wdata     ), 
   .bpf_soc_pcie_slv_wstrb     (bpf_soc_pcie_slv_if.wstrb     ), 
   .bpf_soc_pcie_slv_wvalid    (bpf_soc_pcie_slv_if.wvalid    ), 
   .bpf_soc_pcie_slv_wready    (bpf_soc_pcie_slv_if.wready    ), 
   .bpf_soc_pcie_slv_bresp     (bpf_soc_pcie_slv_if.bresp     ), 
   .bpf_soc_pcie_slv_bvalid    (bpf_soc_pcie_slv_if.bvalid    ), 
   .bpf_soc_pcie_slv_bready    (bpf_soc_pcie_slv_if.bready    ), 
   .bpf_soc_pcie_slv_araddr    (bpf_soc_pcie_slv_if.araddr    ), 
   .bpf_soc_pcie_slv_arprot    (bpf_soc_pcie_slv_if.arprot    ), 
   .bpf_soc_pcie_slv_arvalid   (bpf_soc_pcie_slv_if.arvalid   ), 
   .bpf_soc_pcie_slv_arready   (bpf_soc_pcie_slv_if.arready   ), 
   .bpf_soc_pcie_slv_rdata     (bpf_soc_pcie_slv_if.rdata     ), 
   .bpf_soc_pcie_slv_rresp     (bpf_soc_pcie_slv_if.rresp     ), 
   .bpf_soc_pcie_slv_rvalid    (bpf_soc_pcie_slv_if.rvalid    ), 
   .bpf_soc_pcie_slv_rready    (bpf_soc_pcie_slv_if.rready    ),
 
   .bpf_soc_apf_slv_awaddr    (bpf_soc_apf_slv_if.awaddr     ),
   .bpf_soc_apf_slv_awprot    (bpf_soc_apf_slv_if.awprot     ),
   .bpf_soc_apf_slv_awvalid   (bpf_soc_apf_slv_if.awvalid    ),
   .bpf_soc_apf_slv_awready   (bpf_soc_apf_slv_if.awready    ),
   .bpf_soc_apf_slv_wdata     (bpf_soc_apf_slv_if.wdata      ),
   .bpf_soc_apf_slv_wstrb     (bpf_soc_apf_slv_if.wstrb      ),
   .bpf_soc_apf_slv_wvalid    (bpf_soc_apf_slv_if.wvalid     ),
   .bpf_soc_apf_slv_wready    (bpf_soc_apf_slv_if.wready     ),
   .bpf_soc_apf_slv_bresp     (bpf_soc_apf_slv_if.bresp      ),
   .bpf_soc_apf_slv_bvalid    (bpf_soc_apf_slv_if.bvalid     ),
   .bpf_soc_apf_slv_bready    (bpf_soc_apf_slv_if.bready     ),
   .bpf_soc_apf_slv_araddr    (bpf_soc_apf_slv_if.araddr     ),
   .bpf_soc_apf_slv_arprot    (bpf_soc_apf_slv_if.arprot     ),
   .bpf_soc_apf_slv_arvalid   (bpf_soc_apf_slv_if.arvalid    ),
   .bpf_soc_apf_slv_arready   (bpf_soc_apf_slv_if.arready    ),
   .bpf_soc_apf_slv_rdata     (bpf_soc_apf_slv_if.rdata      ),
   .bpf_soc_apf_slv_rresp     (bpf_soc_apf_slv_if.rresp      ),
   .bpf_soc_apf_slv_rvalid    (bpf_soc_apf_slv_if.rvalid     ),
   .bpf_soc_apf_slv_rready    (bpf_soc_apf_slv_if.rready     ),
   
   .bpf_fme_slv_awaddr        (bpf_fme_slv_if.awaddr     ),
   .bpf_fme_slv_awprot        (bpf_fme_slv_if.awprot     ),
   .bpf_fme_slv_awvalid       (bpf_fme_slv_if.awvalid    ),
   .bpf_fme_slv_awready       (bpf_fme_slv_if.awready    ),
   .bpf_fme_slv_wdata         (bpf_fme_slv_if.wdata      ),
   .bpf_fme_slv_wstrb         (bpf_fme_slv_if.wstrb      ),
   .bpf_fme_slv_wvalid        (bpf_fme_slv_if.wvalid     ),
   .bpf_fme_slv_wready        (bpf_fme_slv_if.wready     ),
   .bpf_fme_slv_bresp         (bpf_fme_slv_if.bresp      ),
   .bpf_fme_slv_bvalid        (bpf_fme_slv_if.bvalid     ),
   .bpf_fme_slv_bready        (bpf_fme_slv_if.bready     ),
   .bpf_fme_slv_araddr        (bpf_fme_slv_if.araddr     ),
   .bpf_fme_slv_arprot        (bpf_fme_slv_if.arprot     ),
   .bpf_fme_slv_arvalid       (bpf_fme_slv_if.arvalid    ),
   .bpf_fme_slv_arready       (bpf_fme_slv_if.arready    ),
   .bpf_fme_slv_rdata         (bpf_fme_slv_if.rdata      ),
   .bpf_fme_slv_rresp         (bpf_fme_slv_if.rresp      ),
   .bpf_fme_slv_rvalid        (bpf_fme_slv_if.rvalid     ),
   .bpf_fme_slv_rready        (bpf_fme_slv_if.rready     ),
    
   .bpf_fme_mst_awaddr        (bpf_fme_mst_if.awaddr     ),
   .bpf_fme_mst_awprot        (bpf_fme_mst_if.awprot     ),
   .bpf_fme_mst_awvalid       (bpf_fme_mst_if.awvalid    ),
   .bpf_fme_mst_awready       (bpf_fme_mst_if.awready    ),
   .bpf_fme_mst_wdata         (bpf_fme_mst_if.wdata      ),
   .bpf_fme_mst_wstrb         (bpf_fme_mst_if.wstrb      ),
   .bpf_fme_mst_wvalid        (bpf_fme_mst_if.wvalid     ),
   .bpf_fme_mst_wready        (bpf_fme_mst_if.wready     ),
   .bpf_fme_mst_bresp         (bpf_fme_mst_if.bresp      ),
   .bpf_fme_mst_bvalid        (bpf_fme_mst_if.bvalid     ),
   .bpf_fme_mst_bready        (bpf_fme_mst_if.bready     ),
   .bpf_fme_mst_araddr        (bpf_fme_mst_if.araddr     ),
   .bpf_fme_mst_arprot        (bpf_fme_mst_if.arprot     ),
   .bpf_fme_mst_arvalid       (bpf_fme_mst_if.arvalid    ),
   .bpf_fme_mst_arready       (bpf_fme_mst_if.arready    ),
   .bpf_fme_mst_rdata         (bpf_fme_mst_if.rdata      ),
   .bpf_fme_mst_rresp         (bpf_fme_mst_if.rresp      ),
   .bpf_fme_mst_rvalid        (bpf_fme_mst_if.rvalid     ),
   .bpf_fme_mst_rready        (bpf_fme_mst_if.rready     ),

   .bpf_pmci_mst_awaddr        (bpf_pmci_mst_if.awaddr     ),
   .bpf_pmci_mst_awprot        (bpf_pmci_mst_if.awprot     ),
   .bpf_pmci_mst_awvalid       (bpf_pmci_mst_if.awvalid    ),
   .bpf_pmci_mst_awready       (bpf_pmci_mst_if.awready    ),
   .bpf_pmci_mst_wdata         (bpf_pmci_mst_if.wdata      ),
   .bpf_pmci_mst_wstrb         (bpf_pmci_mst_if.wstrb      ),
   .bpf_pmci_mst_wvalid        (bpf_pmci_mst_if.wvalid     ),
   .bpf_pmci_mst_wready        (bpf_pmci_mst_if.wready     ),
   .bpf_pmci_mst_bresp         (bpf_pmci_mst_if.bresp      ),
   .bpf_pmci_mst_bvalid        (bpf_pmci_mst_if.bvalid     ),
   .bpf_pmci_mst_bready        (bpf_pmci_mst_if.bready     ),
   .bpf_pmci_mst_araddr        (bpf_pmci_mst_if.araddr     ),
   .bpf_pmci_mst_arprot        (bpf_pmci_mst_if.arprot     ),
   .bpf_pmci_mst_arvalid       (bpf_pmci_mst_if.arvalid    ),
   .bpf_pmci_mst_arready       (bpf_pmci_mst_if.arready    ),
   .bpf_pmci_mst_rdata         (bpf_pmci_mst_if.rdata      ),
   .bpf_pmci_mst_rresp         (bpf_pmci_mst_if.rresp      ),
   .bpf_pmci_mst_rvalid        (bpf_pmci_mst_if.rvalid     ),
   .bpf_pmci_mst_rready        (bpf_pmci_mst_if.rready     ),

   
   .bpf_hssi_slv_awaddr       (bpf_hssi_slv_if.awaddr     ),
   .bpf_hssi_slv_awprot       (bpf_hssi_slv_if.awprot     ),
   .bpf_hssi_slv_awvalid      (bpf_hssi_slv_if.awvalid    ),
   .bpf_hssi_slv_awready      (bpf_hssi_slv_if.awready    ),
   .bpf_hssi_slv_wdata        (bpf_hssi_slv_if.wdata      ),
   .bpf_hssi_slv_wstrb        (bpf_hssi_slv_if.wstrb      ),
   .bpf_hssi_slv_wvalid       (bpf_hssi_slv_if.wvalid     ),
   .bpf_hssi_slv_wready       (bpf_hssi_slv_if.wready     ),
   .bpf_hssi_slv_bresp        (bpf_hssi_slv_if.bresp      ),
   .bpf_hssi_slv_bvalid       (bpf_hssi_slv_if.bvalid     ),
   .bpf_hssi_slv_bready       (bpf_hssi_slv_if.bready     ),
   .bpf_hssi_slv_araddr       (bpf_hssi_slv_if.araddr     ),
   .bpf_hssi_slv_arprot       (bpf_hssi_slv_if.arprot     ),
   .bpf_hssi_slv_arvalid      (bpf_hssi_slv_if.arvalid    ),
   .bpf_hssi_slv_arready      (bpf_hssi_slv_if.arready    ),
   .bpf_hssi_slv_rdata        (bpf_hssi_slv_if.rdata      ),
   .bpf_hssi_slv_rresp        (bpf_hssi_slv_if.rresp      ),
   .bpf_hssi_slv_rvalid       (bpf_hssi_slv_if.rvalid     ),
   .bpf_hssi_slv_rready       (bpf_hssi_slv_if.rready     ),
 
   .bpf_qsfp0_slv_awaddr       (bpf_qsfp0_slv_if.awaddr     ),
   .bpf_qsfp0_slv_awprot       (bpf_qsfp0_slv_if.awprot     ),
   .bpf_qsfp0_slv_awvalid      (bpf_qsfp0_slv_if.awvalid    ),
   .bpf_qsfp0_slv_awready      (bpf_qsfp0_slv_if.awready    ),
   .bpf_qsfp0_slv_wdata        (bpf_qsfp0_slv_if.wdata      ),
   .bpf_qsfp0_slv_wstrb        (bpf_qsfp0_slv_if.wstrb      ),
   .bpf_qsfp0_slv_wvalid       (bpf_qsfp0_slv_if.wvalid     ),
   .bpf_qsfp0_slv_wready       (bpf_qsfp0_slv_if.wready     ),
   .bpf_qsfp0_slv_bresp        (bpf_qsfp0_slv_if.bresp      ),
   .bpf_qsfp0_slv_bvalid       (bpf_qsfp0_slv_if.bvalid     ),
   .bpf_qsfp0_slv_bready       (bpf_qsfp0_slv_if.bready     ),
   .bpf_qsfp0_slv_araddr       (bpf_qsfp0_slv_if.araddr     ),
   .bpf_qsfp0_slv_arprot       (bpf_qsfp0_slv_if.arprot     ),
   .bpf_qsfp0_slv_arvalid      (bpf_qsfp0_slv_if.arvalid    ),
   .bpf_qsfp0_slv_arready      (bpf_qsfp0_slv_if.arready    ),
   .bpf_qsfp0_slv_rdata        (bpf_qsfp0_slv_if.rdata      ),
   .bpf_qsfp0_slv_rresp        (bpf_qsfp0_slv_if.rresp      ),
   .bpf_qsfp0_slv_rvalid       (bpf_qsfp0_slv_if.rvalid     ),
   .bpf_qsfp0_slv_rready       (bpf_qsfp0_slv_if.rready     ),
 
   .bpf_qsfp1_slv_awaddr       (bpf_qsfp1_slv_if.awaddr     ),
   .bpf_qsfp1_slv_awprot       (bpf_qsfp1_slv_if.awprot     ),
   .bpf_qsfp1_slv_awvalid      (bpf_qsfp1_slv_if.awvalid    ),
   .bpf_qsfp1_slv_awready      (bpf_qsfp1_slv_if.awready    ),
   .bpf_qsfp1_slv_wdata        (bpf_qsfp1_slv_if.wdata      ),
   .bpf_qsfp1_slv_wstrb        (bpf_qsfp1_slv_if.wstrb      ),
   .bpf_qsfp1_slv_wvalid       (bpf_qsfp1_slv_if.wvalid     ),
   .bpf_qsfp1_slv_wready       (bpf_qsfp1_slv_if.wready     ),
   .bpf_qsfp1_slv_bresp        (bpf_qsfp1_slv_if.bresp      ),
   .bpf_qsfp1_slv_bvalid       (bpf_qsfp1_slv_if.bvalid     ),
   .bpf_qsfp1_slv_bready       (bpf_qsfp1_slv_if.bready     ),
   .bpf_qsfp1_slv_araddr       (bpf_qsfp1_slv_if.araddr     ),
   .bpf_qsfp1_slv_arprot       (bpf_qsfp1_slv_if.arprot     ),
   .bpf_qsfp1_slv_arvalid      (bpf_qsfp1_slv_if.arvalid    ),
   .bpf_qsfp1_slv_arready      (bpf_qsfp1_slv_if.arready    ),
   .bpf_qsfp1_slv_rdata        (bpf_qsfp1_slv_if.rdata      ),
   .bpf_qsfp1_slv_rresp        (bpf_qsfp1_slv_if.rresp      ),
   .bpf_qsfp1_slv_rvalid       (bpf_qsfp1_slv_if.rvalid     ),
   .bpf_qsfp1_slv_rready       (bpf_qsfp1_slv_if.rready     ),

   .bpf_emif_slv_awaddr    (bpf_emif_slv_if.awaddr    ), 
   .bpf_emif_slv_awprot    (bpf_emif_slv_if.awprot    ), 
   .bpf_emif_slv_awvalid   (bpf_emif_slv_if.awvalid   ), 
   .bpf_emif_slv_awready   (bpf_emif_slv_if.awready   ), 
   .bpf_emif_slv_wdata     (bpf_emif_slv_if.wdata     ), 
   .bpf_emif_slv_wstrb     (bpf_emif_slv_if.wstrb     ), 
   .bpf_emif_slv_wvalid    (bpf_emif_slv_if.wvalid    ), 
   .bpf_emif_slv_wready    (bpf_emif_slv_if.wready    ), 
   .bpf_emif_slv_bresp     (bpf_emif_slv_if.bresp     ), 
   .bpf_emif_slv_bvalid    (bpf_emif_slv_if.bvalid    ), 
   .bpf_emif_slv_bready    (bpf_emif_slv_if.bready    ), 
   .bpf_emif_slv_araddr    (bpf_emif_slv_if.araddr    ), 
   .bpf_emif_slv_arprot    (bpf_emif_slv_if.arprot    ), 
   .bpf_emif_slv_arvalid   (bpf_emif_slv_if.arvalid   ), 
   .bpf_emif_slv_arready   (bpf_emif_slv_if.arready   ), 
   .bpf_emif_slv_rdata     (bpf_emif_slv_if.rdata     ), 
   .bpf_emif_slv_rresp     (bpf_emif_slv_if.rresp     ), 
   .bpf_emif_slv_rvalid    (bpf_emif_slv_if.rvalid    ), 
   .bpf_emif_slv_rready    (bpf_emif_slv_if.rready    ),

   .bpf_pmci_slv_awaddr    (bpf_pmci_slv_if.awaddr     ),
   .bpf_pmci_slv_awprot    (bpf_pmci_slv_if.awprot     ),
   .bpf_pmci_slv_awvalid   (bpf_pmci_slv_if.awvalid    ),
   .bpf_pmci_slv_awready   (bpf_pmci_slv_if.awready    ),
   .bpf_pmci_slv_wdata     (bpf_pmci_slv_if.wdata      ),
   .bpf_pmci_slv_wstrb     (bpf_pmci_slv_if.wstrb      ),
   .bpf_pmci_slv_wvalid    (bpf_pmci_slv_if.wvalid     ),
   .bpf_pmci_slv_wready    (bpf_pmci_slv_if.wready     ),
   .bpf_pmci_slv_bresp     (bpf_pmci_slv_if.bresp      ),
   .bpf_pmci_slv_bvalid    (bpf_pmci_slv_if.bvalid     ),
   .bpf_pmci_slv_bready    (bpf_pmci_slv_if.bready     ),
   .bpf_pmci_slv_araddr    (bpf_pmci_slv_if.araddr     ),
   .bpf_pmci_slv_arprot    (bpf_pmci_slv_if.arprot     ),
   .bpf_pmci_slv_arvalid   (bpf_pmci_slv_if.arvalid    ),
   .bpf_pmci_slv_arready   (bpf_pmci_slv_if.arready    ),
   .bpf_pmci_slv_rdata     (bpf_pmci_slv_if.rdata      ),
   .bpf_pmci_slv_rresp     (bpf_pmci_slv_if.rresp      ),
   .bpf_pmci_slv_rvalid    (bpf_pmci_slv_if.rvalid     ),
   .bpf_pmci_slv_rready    (bpf_pmci_slv_if.rready     ),

   .bpf_host_apf_slv_awaddr    (bpf_host_apf_slv_if.awaddr     ),
   .bpf_host_apf_slv_awprot    (bpf_host_apf_slv_if.awprot     ),
   .bpf_host_apf_slv_awvalid   (bpf_host_apf_slv_if.awvalid    ),
   .bpf_host_apf_slv_awready   (bpf_host_apf_slv_if.awready    ),
   .bpf_host_apf_slv_wdata     (bpf_host_apf_slv_if.wdata      ),
   .bpf_host_apf_slv_wstrb     (bpf_host_apf_slv_if.wstrb      ),
   .bpf_host_apf_slv_wvalid    (bpf_host_apf_slv_if.wvalid     ),
   .bpf_host_apf_slv_wready    (bpf_host_apf_slv_if.wready     ),
   .bpf_host_apf_slv_bresp     (bpf_host_apf_slv_if.bresp      ),
   .bpf_host_apf_slv_bvalid    (bpf_host_apf_slv_if.bvalid     ),
   .bpf_host_apf_slv_bready    (bpf_host_apf_slv_if.bready     ),
   .bpf_host_apf_slv_araddr    (bpf_host_apf_slv_if.araddr     ),
   .bpf_host_apf_slv_arprot    (bpf_host_apf_slv_if.arprot     ),
   .bpf_host_apf_slv_arvalid   (bpf_host_apf_slv_if.arvalid    ),
   .bpf_host_apf_slv_arready   (bpf_host_apf_slv_if.arready    ),
   .bpf_host_apf_slv_rdata     (bpf_host_apf_slv_if.rdata      ),
   .bpf_host_apf_slv_rresp     (bpf_host_apf_slv_if.rresp      ),
   .bpf_host_apf_slv_rvalid    (bpf_host_apf_slv_if.rvalid     ),
   .bpf_host_apf_slv_rready    (bpf_host_apf_slv_if.rready     )

   );

endmodule
